-- VGASubsystem.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity VGASubsystem is
	port (
		char_buffer_control_slave_address    : in  std_logic                     := '0';             -- char_buffer_control_slave.address
		char_buffer_control_slave_byteenable : in  std_logic_vector(3 downto 0)  := (others => '0'); --                          .byteenable
		char_buffer_control_slave_chipselect : in  std_logic                     := '0';             --                          .chipselect
		char_buffer_control_slave_read       : in  std_logic                     := '0';             --                          .read
		char_buffer_control_slave_write      : in  std_logic                     := '0';             --                          .write
		char_buffer_control_slave_writedata  : in  std_logic_vector(31 downto 0) := (others => '0'); --                          .writedata
		char_buffer_control_slave_readdata   : out std_logic_vector(31 downto 0);                    --                          .readdata
		char_buffersource_slave_byteenable   : in  std_logic                     := '0';             --   char_buffersource_slave.byteenable
		char_buffersource_slave_chipselect   : in  std_logic                     := '0';             --                          .chipselect
		char_buffersource_slave_read         : in  std_logic                     := '0';             --                          .read
		char_buffersource_slave_write        : in  std_logic                     := '0';             --                          .write
		char_buffersource_slave_writedata    : in  std_logic_vector(7 downto 0)  := (others => '0'); --                          .writedata
		char_buffersource_slave_readdata     : out std_logic_vector(7 downto 0);                     --                          .readdata
		char_buffersource_slave_waitrequest  : out std_logic;                                        --                          .waitrequest
		char_buffersource_slave_address      : in  std_logic_vector(12 downto 0) := (others => '0'); --                          .address
		pixel_buffer_master_readdatavalid    : in  std_logic                     := '0';             --       pixel_buffer_master.readdatavalid
		pixel_buffer_master_waitrequest      : in  std_logic                     := '0';             --                          .waitrequest
		pixel_buffer_master_address          : out std_logic_vector(31 downto 0);                    --                          .address
		pixel_buffer_master_lock             : out std_logic;                                        --                          .lock
		pixel_buffer_master_read             : out std_logic;                                        --                          .read
		pixel_buffer_master_readdata         : in  std_logic_vector(15 downto 0) := (others => '0'); --                          .readdata
		pixel_buffer_slave_address           : in  std_logic_vector(1 downto 0)  := (others => '0'); --        pixel_buffer_slave.address
		pixel_buffer_slave_byteenable        : in  std_logic_vector(3 downto 0)  := (others => '0'); --                          .byteenable
		pixel_buffer_slave_read              : in  std_logic                     := '0';             --                          .read
		pixel_buffer_slave_write             : in  std_logic                     := '0';             --                          .write
		pixel_buffer_slave_writedata         : in  std_logic_vector(31 downto 0) := (others => '0'); --                          .writedata
		pixel_buffer_slave_readdata          : out std_logic_vector(31 downto 0);                    --                          .readdata
		rgb_resampler_slave_read             : in  std_logic                     := '0';             --       rgb_resampler_slave.read
		rgb_resampler_slave_readdata         : out std_logic_vector(31 downto 0);                    --                          .readdata
		sys_clk_clk                          : in  std_logic                     := '0';             --                   sys_clk.clk
		sys_reset_reset_n                    : in  std_logic                     := '0';             --                 sys_reset.reset_n
		vga_CLK                              : out std_logic;                                        --                       vga.CLK
		vga_HS                               : out std_logic;                                        --                          .HS
		vga_VS                               : out std_logic;                                        --                          .VS
		vga_BLANK                            : out std_logic;                                        --                          .BLANK
		vga_SYNC                             : out std_logic;                                        --                          .SYNC
		vga_R                                : out std_logic_vector(7 downto 0);                     --                          .R
		vga_G                                : out std_logic_vector(7 downto 0);                     --                          .G
		vga_B                                : out std_logic_vector(7 downto 0);                     --                          .B
		vga_clk_clk                          : in  std_logic                     := '0';             --                   vga_clk.clk
		vga_reset_reset_n                    : in  std_logic                     := '0'              --                 vga_reset.reset_n
	);
end entity VGASubsystem;

architecture rtl of VGASubsystem is
	component VGASubsystem_Alpha_Blender is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			foreground_data          : in  std_logic_vector(39 downto 0) := (others => 'X'); -- data
			foreground_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			foreground_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			foreground_valid         : in  std_logic                     := 'X';             -- valid
			foreground_ready         : out std_logic;                                        -- ready
			background_data          : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			background_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			background_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			background_valid         : in  std_logic                     := 'X';             -- valid
			background_ready         : out std_logic;                                        -- ready
			output_ready             : in  std_logic                     := 'X';             -- ready
			output_data              : out std_logic_vector(29 downto 0);                    -- data
			output_startofpacket     : out std_logic;                                        -- startofpacket
			output_endofpacket       : out std_logic;                                        -- endofpacket
			output_valid             : out std_logic                                         -- valid
		);
	end component VGASubsystem_Alpha_Blender;

	component VGASubsystem_Character_Buffer is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			ctrl_address         : in  std_logic                     := 'X';             -- address
			ctrl_byteenable      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			ctrl_chipselect      : in  std_logic                     := 'X';             -- chipselect
			ctrl_read            : in  std_logic                     := 'X';             -- read
			ctrl_write           : in  std_logic                     := 'X';             -- write
			ctrl_writedata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			ctrl_readdata        : out std_logic_vector(31 downto 0);                    -- readdata
			buf_byteenable       : in  std_logic                     := 'X';             -- byteenable
			buf_chipselect       : in  std_logic                     := 'X';             -- chipselect
			buf_read             : in  std_logic                     := 'X';             -- read
			buf_write            : in  std_logic                     := 'X';             -- write
			buf_writedata        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			buf_readdata         : out std_logic_vector(7 downto 0);                     -- readdata
			buf_waitrequest      : out std_logic;                                        -- waitrequest
			buf_address          : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			stream_ready         : in  std_logic                     := 'X';             -- ready
			stream_startofpacket : out std_logic;                                        -- startofpacket
			stream_endofpacket   : out std_logic;                                        -- endofpacket
			stream_valid         : out std_logic;                                        -- valid
			stream_data          : out std_logic_vector(39 downto 0)                     -- data
		);
	end component VGASubsystem_Character_Buffer;

	component VGASubsystem_Dual_Clock_FIFO is
		port (
			clk_stream_in            : in  std_logic                     := 'X';             -- clk
			reset_stream_in          : in  std_logic                     := 'X';             -- reset
			clk_stream_out           : in  std_logic                     := 'X';             -- clk
			reset_stream_out         : in  std_logic                     := 'X';             -- reset
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_data           : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(29 downto 0)                     -- data
		);
	end component VGASubsystem_Dual_Clock_FIFO;

	component VGASubsystem_Pixel_Buffer is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_arbiterlock   : out std_logic;                                        -- lock
			master_read          : out std_logic;                                        -- read
			master_readdata      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			slave_address        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			slave_byteenable     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			slave_read           : in  std_logic                     := 'X';             -- read
			slave_write          : in  std_logic                     := 'X';             -- write
			slave_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			stream_ready         : in  std_logic                     := 'X';             -- ready
			stream_startofpacket : out std_logic;                                        -- startofpacket
			stream_endofpacket   : out std_logic;                                        -- endofpacket
			stream_valid         : out std_logic;                                        -- valid
			stream_data          : out std_logic_vector(15 downto 0)                     -- data
		);
	end component VGASubsystem_Pixel_Buffer;

	component VGASubsystem_Resampler is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_data           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			slave_read               : in  std_logic                     := 'X';             -- read
			slave_readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(29 downto 0)                     -- data
		);
	end component VGASubsystem_Resampler;

	component VGASubsystem_VGA_Controller is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X';             -- reset
			data          : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			startofpacket : in  std_logic                     := 'X';             -- startofpacket
			endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			valid         : in  std_logic                     := 'X';             -- valid
			ready         : out std_logic;                                        -- ready
			VGA_CLK       : out std_logic;                                        -- export
			VGA_HS        : out std_logic;                                        -- export
			VGA_VS        : out std_logic;                                        -- export
			VGA_BLANK     : out std_logic;                                        -- export
			VGA_SYNC      : out std_logic;                                        -- export
			VGA_R         : out std_logic_vector(7 downto 0);                     -- export
			VGA_G         : out std_logic_vector(7 downto 0);                     -- export
			VGA_B         : out std_logic_vector(7 downto 0)                      -- export
		);
	end component VGASubsystem_VGA_Controller;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal alpha_blender_avalon_blended_source_valid             : std_logic;                     -- Alpha_Blender:output_valid -> Dual_Clock_FIFO:stream_in_valid
	signal alpha_blender_avalon_blended_source_data              : std_logic_vector(29 downto 0); -- Alpha_Blender:output_data -> Dual_Clock_FIFO:stream_in_data
	signal alpha_blender_avalon_blended_source_ready             : std_logic;                     -- Dual_Clock_FIFO:stream_in_ready -> Alpha_Blender:output_ready
	signal alpha_blender_avalon_blended_source_startofpacket     : std_logic;                     -- Alpha_Blender:output_startofpacket -> Dual_Clock_FIFO:stream_in_startofpacket
	signal alpha_blender_avalon_blended_source_endofpacket       : std_logic;                     -- Alpha_Blender:output_endofpacket -> Dual_Clock_FIFO:stream_in_endofpacket
	signal character_buffer_avalon_char_source_valid             : std_logic;                     -- Character_Buffer:stream_valid -> Alpha_Blender:foreground_valid
	signal character_buffer_avalon_char_source_data              : std_logic_vector(39 downto 0); -- Character_Buffer:stream_data -> Alpha_Blender:foreground_data
	signal character_buffer_avalon_char_source_ready             : std_logic;                     -- Alpha_Blender:foreground_ready -> Character_Buffer:stream_ready
	signal character_buffer_avalon_char_source_startofpacket     : std_logic;                     -- Character_Buffer:stream_startofpacket -> Alpha_Blender:foreground_startofpacket
	signal character_buffer_avalon_char_source_endofpacket       : std_logic;                     -- Character_Buffer:stream_endofpacket -> Alpha_Blender:foreground_endofpacket
	signal dual_clock_fifo_avalon_dc_buffer_source_valid         : std_logic;                     -- Dual_Clock_FIFO:stream_out_valid -> VGA_Controller:valid
	signal dual_clock_fifo_avalon_dc_buffer_source_data          : std_logic_vector(29 downto 0); -- Dual_Clock_FIFO:stream_out_data -> VGA_Controller:data
	signal dual_clock_fifo_avalon_dc_buffer_source_ready         : std_logic;                     -- VGA_Controller:ready -> Dual_Clock_FIFO:stream_out_ready
	signal dual_clock_fifo_avalon_dc_buffer_source_startofpacket : std_logic;                     -- Dual_Clock_FIFO:stream_out_startofpacket -> VGA_Controller:startofpacket
	signal dual_clock_fifo_avalon_dc_buffer_source_endofpacket   : std_logic;                     -- Dual_Clock_FIFO:stream_out_endofpacket -> VGA_Controller:endofpacket
	signal pixel_buffer_avalon_pixel_source_valid                : std_logic;                     -- Pixel_Buffer:stream_valid -> Resampler:stream_in_valid
	signal pixel_buffer_avalon_pixel_source_data                 : std_logic_vector(15 downto 0); -- Pixel_Buffer:stream_data -> Resampler:stream_in_data
	signal pixel_buffer_avalon_pixel_source_ready                : std_logic;                     -- Resampler:stream_in_ready -> Pixel_Buffer:stream_ready
	signal pixel_buffer_avalon_pixel_source_startofpacket        : std_logic;                     -- Pixel_Buffer:stream_startofpacket -> Resampler:stream_in_startofpacket
	signal pixel_buffer_avalon_pixel_source_endofpacket          : std_logic;                     -- Pixel_Buffer:stream_endofpacket -> Resampler:stream_in_endofpacket
	signal resampler_avalon_rgb_source_valid                     : std_logic;                     -- Resampler:stream_out_valid -> Alpha_Blender:background_valid
	signal resampler_avalon_rgb_source_data                      : std_logic_vector(29 downto 0); -- Resampler:stream_out_data -> Alpha_Blender:background_data
	signal resampler_avalon_rgb_source_ready                     : std_logic;                     -- Alpha_Blender:background_ready -> Resampler:stream_out_ready
	signal resampler_avalon_rgb_source_startofpacket             : std_logic;                     -- Resampler:stream_out_startofpacket -> Alpha_Blender:background_startofpacket
	signal resampler_avalon_rgb_source_endofpacket               : std_logic;                     -- Resampler:stream_out_endofpacket -> Alpha_Blender:background_endofpacket
	signal rst_controller_reset_out_reset                        : std_logic;                     -- rst_controller:reset_out -> [Alpha_Blender:reset, Character_Buffer:reset, Dual_Clock_FIFO:reset_stream_in, Pixel_Buffer:reset, Resampler:reset]
	signal rst_controller_001_reset_out_reset                    : std_logic;                     -- rst_controller_001:reset_out -> [Dual_Clock_FIFO:reset_stream_out, VGA_Controller:reset]
	signal sys_reset_reset_n_ports_inv                           : std_logic;                     -- sys_reset_reset_n:inv -> rst_controller:reset_in0
	signal vga_reset_reset_n_ports_inv                           : std_logic;                     -- vga_reset_reset_n:inv -> rst_controller_001:reset_in0

begin

	alpha_blender : component VGASubsystem_Alpha_Blender
		port map (
			clk                      => sys_clk_clk,                                       --                    clk.clk
			reset                    => rst_controller_reset_out_reset,                    --                  reset.reset
			foreground_data          => character_buffer_avalon_char_source_data,          -- avalon_foreground_sink.data
			foreground_startofpacket => character_buffer_avalon_char_source_startofpacket, --                       .startofpacket
			foreground_endofpacket   => character_buffer_avalon_char_source_endofpacket,   --                       .endofpacket
			foreground_valid         => character_buffer_avalon_char_source_valid,         --                       .valid
			foreground_ready         => character_buffer_avalon_char_source_ready,         --                       .ready
			background_data          => resampler_avalon_rgb_source_data,                  -- avalon_background_sink.data
			background_startofpacket => resampler_avalon_rgb_source_startofpacket,         --                       .startofpacket
			background_endofpacket   => resampler_avalon_rgb_source_endofpacket,           --                       .endofpacket
			background_valid         => resampler_avalon_rgb_source_valid,                 --                       .valid
			background_ready         => resampler_avalon_rgb_source_ready,                 --                       .ready
			output_ready             => alpha_blender_avalon_blended_source_ready,         --  avalon_blended_source.ready
			output_data              => alpha_blender_avalon_blended_source_data,          --                       .data
			output_startofpacket     => alpha_blender_avalon_blended_source_startofpacket, --                       .startofpacket
			output_endofpacket       => alpha_blender_avalon_blended_source_endofpacket,   --                       .endofpacket
			output_valid             => alpha_blender_avalon_blended_source_valid          --                       .valid
		);

	character_buffer : component VGASubsystem_Character_Buffer
		port map (
			clk                  => sys_clk_clk,                                       --                       clk.clk
			reset                => rst_controller_reset_out_reset,                    --                     reset.reset
			ctrl_address         => char_buffer_control_slave_address,                 -- avalon_char_control_slave.address
			ctrl_byteenable      => char_buffer_control_slave_byteenable,              --                          .byteenable
			ctrl_chipselect      => char_buffer_control_slave_chipselect,              --                          .chipselect
			ctrl_read            => char_buffer_control_slave_read,                    --                          .read
			ctrl_write           => char_buffer_control_slave_write,                   --                          .write
			ctrl_writedata       => char_buffer_control_slave_writedata,               --                          .writedata
			ctrl_readdata        => char_buffer_control_slave_readdata,                --                          .readdata
			buf_byteenable       => char_buffersource_slave_byteenable,                --  avalon_char_buffer_slave.byteenable
			buf_chipselect       => char_buffersource_slave_chipselect,                --                          .chipselect
			buf_read             => char_buffersource_slave_read,                      --                          .read
			buf_write            => char_buffersource_slave_write,                     --                          .write
			buf_writedata        => char_buffersource_slave_writedata,                 --                          .writedata
			buf_readdata         => char_buffersource_slave_readdata,                  --                          .readdata
			buf_waitrequest      => char_buffersource_slave_waitrequest,               --                          .waitrequest
			buf_address          => char_buffersource_slave_address,                   --                          .address
			stream_ready         => character_buffer_avalon_char_source_ready,         --        avalon_char_source.ready
			stream_startofpacket => character_buffer_avalon_char_source_startofpacket, --                          .startofpacket
			stream_endofpacket   => character_buffer_avalon_char_source_endofpacket,   --                          .endofpacket
			stream_valid         => character_buffer_avalon_char_source_valid,         --                          .valid
			stream_data          => character_buffer_avalon_char_source_data           --                          .data
		);

	dual_clock_fifo : component VGASubsystem_Dual_Clock_FIFO
		port map (
			clk_stream_in            => sys_clk_clk,                                           --         clock_stream_in.clk
			reset_stream_in          => rst_controller_reset_out_reset,                        --         reset_stream_in.reset
			clk_stream_out           => vga_clk_clk,                                           --        clock_stream_out.clk
			reset_stream_out         => rst_controller_001_reset_out_reset,                    --        reset_stream_out.reset
			stream_in_ready          => alpha_blender_avalon_blended_source_ready,             --   avalon_dc_buffer_sink.ready
			stream_in_startofpacket  => alpha_blender_avalon_blended_source_startofpacket,     --                        .startofpacket
			stream_in_endofpacket    => alpha_blender_avalon_blended_source_endofpacket,       --                        .endofpacket
			stream_in_valid          => alpha_blender_avalon_blended_source_valid,             --                        .valid
			stream_in_data           => alpha_blender_avalon_blended_source_data,              --                        .data
			stream_out_ready         => dual_clock_fifo_avalon_dc_buffer_source_ready,         -- avalon_dc_buffer_source.ready
			stream_out_startofpacket => dual_clock_fifo_avalon_dc_buffer_source_startofpacket, --                        .startofpacket
			stream_out_endofpacket   => dual_clock_fifo_avalon_dc_buffer_source_endofpacket,   --                        .endofpacket
			stream_out_valid         => dual_clock_fifo_avalon_dc_buffer_source_valid,         --                        .valid
			stream_out_data          => dual_clock_fifo_avalon_dc_buffer_source_data           --                        .data
		);

	pixel_buffer : component VGASubsystem_Pixel_Buffer
		port map (
			clk                  => sys_clk_clk,                                    --                     clk.clk
			reset                => rst_controller_reset_out_reset,                 --                   reset.reset
			master_readdatavalid => pixel_buffer_master_readdatavalid,              -- avalon_pixel_dma_master.readdatavalid
			master_waitrequest   => pixel_buffer_master_waitrequest,                --                        .waitrequest
			master_address       => pixel_buffer_master_address,                    --                        .address
			master_arbiterlock   => pixel_buffer_master_lock,                       --                        .lock
			master_read          => pixel_buffer_master_read,                       --                        .read
			master_readdata      => pixel_buffer_master_readdata,                   --                        .readdata
			slave_address        => pixel_buffer_slave_address,                     --    avalon_control_slave.address
			slave_byteenable     => pixel_buffer_slave_byteenable,                  --                        .byteenable
			slave_read           => pixel_buffer_slave_read,                        --                        .read
			slave_write          => pixel_buffer_slave_write,                       --                        .write
			slave_writedata      => pixel_buffer_slave_writedata,                   --                        .writedata
			slave_readdata       => pixel_buffer_slave_readdata,                    --                        .readdata
			stream_ready         => pixel_buffer_avalon_pixel_source_ready,         --     avalon_pixel_source.ready
			stream_startofpacket => pixel_buffer_avalon_pixel_source_startofpacket, --                        .startofpacket
			stream_endofpacket   => pixel_buffer_avalon_pixel_source_endofpacket,   --                        .endofpacket
			stream_valid         => pixel_buffer_avalon_pixel_source_valid,         --                        .valid
			stream_data          => pixel_buffer_avalon_pixel_source_data           --                        .data
		);

	resampler : component VGASubsystem_Resampler
		port map (
			clk                      => sys_clk_clk,                                    --               clk.clk
			reset                    => rst_controller_reset_out_reset,                 --             reset.reset
			stream_in_startofpacket  => pixel_buffer_avalon_pixel_source_startofpacket, --   avalon_rgb_sink.startofpacket
			stream_in_endofpacket    => pixel_buffer_avalon_pixel_source_endofpacket,   --                  .endofpacket
			stream_in_valid          => pixel_buffer_avalon_pixel_source_valid,         --                  .valid
			stream_in_ready          => pixel_buffer_avalon_pixel_source_ready,         --                  .ready
			stream_in_data           => pixel_buffer_avalon_pixel_source_data,          --                  .data
			slave_read               => rgb_resampler_slave_read,                       --  avalon_rgb_slave.read
			slave_readdata           => rgb_resampler_slave_readdata,                   --                  .readdata
			stream_out_ready         => resampler_avalon_rgb_source_ready,              -- avalon_rgb_source.ready
			stream_out_startofpacket => resampler_avalon_rgb_source_startofpacket,      --                  .startofpacket
			stream_out_endofpacket   => resampler_avalon_rgb_source_endofpacket,        --                  .endofpacket
			stream_out_valid         => resampler_avalon_rgb_source_valid,              --                  .valid
			stream_out_data          => resampler_avalon_rgb_source_data                --                  .data
		);

	vga_controller : component VGASubsystem_VGA_Controller
		port map (
			clk           => vga_clk_clk,                                           --                clk.clk
			reset         => rst_controller_001_reset_out_reset,                    --              reset.reset
			data          => dual_clock_fifo_avalon_dc_buffer_source_data,          --    avalon_vga_sink.data
			startofpacket => dual_clock_fifo_avalon_dc_buffer_source_startofpacket, --                   .startofpacket
			endofpacket   => dual_clock_fifo_avalon_dc_buffer_source_endofpacket,   --                   .endofpacket
			valid         => dual_clock_fifo_avalon_dc_buffer_source_valid,         --                   .valid
			ready         => dual_clock_fifo_avalon_dc_buffer_source_ready,         --                   .ready
			VGA_CLK       => vga_CLK,                                               -- external_interface.export
			VGA_HS        => vga_HS,                                                --                   .export
			VGA_VS        => vga_VS,                                                --                   .export
			VGA_BLANK     => vga_BLANK,                                             --                   .export
			VGA_SYNC      => vga_SYNC,                                              --                   .export
			VGA_R         => vga_R,                                                 --                   .export
			VGA_G         => vga_G,                                                 --                   .export
			VGA_B         => vga_B                                                  --                   .export
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => sys_reset_reset_n_ports_inv,    -- reset_in0.reset
			clk            => sys_clk_clk,                    --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => vga_reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => vga_clk_clk,                        --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	sys_reset_reset_n_ports_inv <= not sys_reset_reset_n;

	vga_reset_reset_n_ports_inv <= not vga_reset_reset_n;

end architecture rtl; -- of VGASubsystem
