-- EV19_SoC.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity EV19_SoC is
	port (
		adc_0_external_interface_sclk : out   std_logic;                                        -- adc_0_external_interface.sclk
		adc_0_external_interface_cs_n : out   std_logic;                                        --                         .cs_n
		adc_0_external_interface_dout : in    std_logic                     := '0';             --                         .dout
		adc_0_external_interface_din  : out   std_logic;                                        --                         .din
		clk_clk                       : in    std_logic                     := '0';             --                      clk.clk
		dip_export                    : in    std_logic_vector(3 downto 0)  := (others => '0'); --                      dip.export
		enablepredictor_config        : in    std_logic                     := '0';             --          enablepredictor.config
		key_export                    : in    std_logic                     := '0';             --                      key.export
		keyboard_CLK                  : inout std_logic                     := '0';             --                 keyboard.CLK
		keyboard_DAT                  : inout std_logic                     := '0';             --                         .DAT
		led_export                    : out   std_logic_vector(7 downto 0);                     --                      led.export
		reset_reset_n                 : in    std_logic                     := '0';             --                    reset.reset_n
		sdram_clk_clk                 : out   std_logic;                                        --                sdram_clk.clk
		sdram_wire_addr               : out   std_logic_vector(12 downto 0);                    --               sdram_wire.addr
		sdram_wire_ba                 : out   std_logic_vector(1 downto 0);                     --                         .ba
		sdram_wire_cas_n              : out   std_logic;                                        --                         .cas_n
		sdram_wire_cke                : out   std_logic;                                        --                         .cke
		sdram_wire_cs_n               : out   std_logic;                                        --                         .cs_n
		sdram_wire_dq                 : inout std_logic_vector(15 downto 0) := (others => '0'); --                         .dq
		sdram_wire_dqm                : out   std_logic_vector(1 downto 0);                     --                         .dqm
		sdram_wire_ras_n              : out   std_logic;                                        --                         .ras_n
		sdram_wire_we_n               : out   std_logic;                                        --                         .we_n
		vga_CLK                       : out   std_logic;                                        --                      vga.CLK
		vga_HS                        : out   std_logic;                                        --                         .HS
		vga_VS                        : out   std_logic;                                        --                         .VS
		vga_BLANK                     : out   std_logic;                                        --                         .BLANK
		vga_SYNC                      : out   std_logic;                                        --                         .SYNC
		vga_R                         : out   std_logic_vector(7 downto 0);                     --                         .R
		vga_G                         : out   std_logic_vector(7 downto 0);                     --                         .G
		vga_B                         : out   std_logic_vector(7 downto 0)                      --                         .B
	);
end entity EV19_SoC;

architecture rtl of EV19_SoC is
	component EV19_SoC_ADC is
		generic (
			board          : string  := "DE10-Standard";
			board_rev      : string  := "Autodetect";
			tsclk          : integer := 0;
			numch          : integer := 0;
			max10pllmultby : integer := 0;
			max10plldivby  : integer := 0
		);
		port (
			clock       : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			address     : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			waitrequest : out std_logic;                                        -- waitrequest
			read        : in  std_logic                     := 'X';             -- read
			adc_sclk    : out std_logic;                                        -- export
			adc_cs_n    : out std_logic;                                        -- export
			adc_dout    : in  std_logic                     := 'X';             -- export
			adc_din     : out std_logic                                         -- export
		);
	end component EV19_SoC_ADC;

	component EV19_SoC_Dip_Switch is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component EV19_SoC_Dip_Switch;

	component Core is
		port (
			reset             : in  std_logic                     := 'X';             -- reset
			dataMemAddress    : out std_logic_vector(31 downto 0);                    -- address
			dataMemByteEnable : out std_logic_vector(3 downto 0);                     -- byteenable
			dataMemReadData   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			dataMemReadReq    : out std_logic;                                        -- read
			dataMemWaitReq    : in  std_logic                     := 'X';             -- waitrequest
			dataMemWriteData  : out std_logic_vector(31 downto 0);                    -- writedata
			dataMemWriteReq   : out std_logic;                                        -- write
			instMemWaitReq    : in  std_logic                     := 'X';             -- waitrequest
			instMemReadData   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			instMemReadReq    : out std_logic;                                        -- read
			instMemByteEnable : out std_logic_vector(3 downto 0);                     -- byteenable
			instMemAddress    : out std_logic_vector(31 downto 0);                    -- address
			clock             : in  std_logic                     := 'X';             -- clk
			enablePredictor   : in  std_logic                     := 'X'              -- config
		);
	end component Core;

	component EV19_SoC_ID is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component EV19_SoC_ID;

	component EV19_SoC_Keyboard is
		port (
			clk         : in    std_logic                     := 'X';             -- clk
			reset       : in    std_logic                     := 'X';             -- reset
			address     : in    std_logic                     := 'X';             -- address
			chipselect  : in    std_logic                     := 'X';             -- chipselect
			byteenable  : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			read        : in    std_logic                     := 'X';             -- read
			write       : in    std_logic                     := 'X';             -- write
			writedata   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata    : out   std_logic_vector(31 downto 0);                    -- readdata
			waitrequest : out   std_logic;                                        -- waitrequest
			irq         : out   std_logic;                                        -- irq
			PS2_CLK     : inout std_logic                     := 'X';             -- export
			PS2_DAT     : inout std_logic                     := 'X'              -- export
		);
	end component EV19_SoC_Keyboard;

	component EV19_SoC_LEDs is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component EV19_SoC_LEDs;

	component EV19_SoC_PLL is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			inclk0             : in  std_logic                     := 'X';             -- clk
			c0                 : out std_logic;                                        -- clk
			c1                 : out std_logic;                                        -- clk
			c2                 : out std_logic;                                        -- clk
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			areset             : in  std_logic                     := 'X';             -- export
			locked             : out std_logic;                                        -- export
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component EV19_SoC_PLL;

	component EV19_SoC_Performance_Counter is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			write         : in  std_logic                     := 'X';             -- write
			writedata     : in  std_logic_vector(31 downto 0) := (others => 'X')  -- writedata
		);
	end component EV19_SoC_Performance_Counter;

	component EV19_SoC_Push_Button is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic                     := 'X'              -- export
		);
	end component EV19_SoC_Push_Button;

	component EV19_SoC_RAM is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component EV19_SoC_RAM;

	component EV19_SoC_ROM is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			address     : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			debugaccess : in  std_logic                     := 'X';             -- debugaccess
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			freeze      : in  std_logic                     := 'X'              -- freeze
		);
	end component EV19_SoC_ROM;

	component EV19_SoC_SDRAM is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(23 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component EV19_SoC_SDRAM;

	component EV19_SoC_Timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component EV19_SoC_Timer;

	component EV19_SoC_VGA is
		port (
			char_buffer_control_slave_address    : in  std_logic                     := 'X';             -- address
			char_buffer_control_slave_byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			char_buffer_control_slave_chipselect : in  std_logic                     := 'X';             -- chipselect
			char_buffer_control_slave_read       : in  std_logic                     := 'X';             -- read
			char_buffer_control_slave_write      : in  std_logic                     := 'X';             -- write
			char_buffer_control_slave_writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			char_buffer_control_slave_readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			char_buffersource_slave_byteenable   : in  std_logic                     := 'X';             -- byteenable
			char_buffersource_slave_chipselect   : in  std_logic                     := 'X';             -- chipselect
			char_buffersource_slave_read         : in  std_logic                     := 'X';             -- read
			char_buffersource_slave_write        : in  std_logic                     := 'X';             -- write
			char_buffersource_slave_writedata    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			char_buffersource_slave_readdata     : out std_logic_vector(7 downto 0);                     -- readdata
			char_buffersource_slave_waitrequest  : out std_logic;                                        -- waitrequest
			char_buffersource_slave_address      : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			pixel_buffer_master_readdatavalid    : in  std_logic                     := 'X';             -- readdatavalid
			pixel_buffer_master_waitrequest      : in  std_logic                     := 'X';             -- waitrequest
			pixel_buffer_master_address          : out std_logic_vector(31 downto 0);                    -- address
			pixel_buffer_master_lock             : out std_logic;                                        -- lock
			pixel_buffer_master_read             : out std_logic;                                        -- read
			pixel_buffer_master_readdata         : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			pixel_buffer_slave_address           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			pixel_buffer_slave_byteenable        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			pixel_buffer_slave_read              : in  std_logic                     := 'X';             -- read
			pixel_buffer_slave_write             : in  std_logic                     := 'X';             -- write
			pixel_buffer_slave_writedata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			pixel_buffer_slave_readdata          : out std_logic_vector(31 downto 0);                    -- readdata
			rgb_resampler_slave_read             : in  std_logic                     := 'X';             -- read
			rgb_resampler_slave_readdata         : out std_logic_vector(31 downto 0);                    -- readdata
			sys_clk_clk                          : in  std_logic                     := 'X';             -- clk
			sys_reset_reset_n                    : in  std_logic                     := 'X';             -- reset_n
			vga_CLK                              : out std_logic;                                        -- CLK
			vga_HS                               : out std_logic;                                        -- HS
			vga_VS                               : out std_logic;                                        -- VS
			vga_BLANK                            : out std_logic;                                        -- BLANK
			vga_SYNC                             : out std_logic;                                        -- SYNC
			vga_R                                : out std_logic_vector(7 downto 0);                     -- R
			vga_G                                : out std_logic_vector(7 downto 0);                     -- G
			vga_B                                : out std_logic_vector(7 downto 0);                     -- B
			vga_clk_clk                          : in  std_logic                     := 'X';             -- clk
			vga_reset_reset_n                    : in  std_logic                     := 'X'              -- reset_n
		);
	end component EV19_SoC_VGA;

	component EV19_SoC_mm_interconnect_0 is
		port (
			PLL_c0_clk                                      : in  std_logic                     := 'X';             -- clk
			EV19_Core_0_reset_reset_bridge_in_reset_reset   : in  std_logic                     := 'X';             -- reset
			VGA_sys_reset_reset_bridge_in_reset_reset       : in  std_logic                     := 'X';             -- reset
			EV19_Core_0_Data_Master_address                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			EV19_Core_0_Data_Master_waitrequest             : out std_logic;                                        -- waitrequest
			EV19_Core_0_Data_Master_byteenable              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			EV19_Core_0_Data_Master_read                    : in  std_logic                     := 'X';             -- read
			EV19_Core_0_Data_Master_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			EV19_Core_0_Data_Master_write                   : in  std_logic                     := 'X';             -- write
			EV19_Core_0_Data_Master_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			EV19_Core_0_Instruction_Master_address          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			EV19_Core_0_Instruction_Master_waitrequest      : out std_logic;                                        -- waitrequest
			EV19_Core_0_Instruction_Master_byteenable       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			EV19_Core_0_Instruction_Master_read             : in  std_logic                     := 'X';             -- read
			EV19_Core_0_Instruction_Master_readdata         : out std_logic_vector(31 downto 0);                    -- readdata
			VGA_pixel_buffer_master_address                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			VGA_pixel_buffer_master_waitrequest             : out std_logic;                                        -- waitrequest
			VGA_pixel_buffer_master_read                    : in  std_logic                     := 'X';             -- read
			VGA_pixel_buffer_master_readdata                : out std_logic_vector(15 downto 0);                    -- readdata
			VGA_pixel_buffer_master_readdatavalid           : out std_logic;                                        -- readdatavalid
			VGA_pixel_buffer_master_lock                    : in  std_logic                     := 'X';             -- lock
			ADC_adc_slave_address                           : out std_logic_vector(2 downto 0);                     -- address
			ADC_adc_slave_write                             : out std_logic;                                        -- write
			ADC_adc_slave_read                              : out std_logic;                                        -- read
			ADC_adc_slave_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ADC_adc_slave_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			ADC_adc_slave_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			Dip_Switch_s1_address                           : out std_logic_vector(1 downto 0);                     -- address
			Dip_Switch_s1_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ID_control_slave_address                        : out std_logic_vector(0 downto 0);                     -- address
			ID_control_slave_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Keyboard_avalon_ps2_slave_address               : out std_logic_vector(0 downto 0);                     -- address
			Keyboard_avalon_ps2_slave_write                 : out std_logic;                                        -- write
			Keyboard_avalon_ps2_slave_read                  : out std_logic;                                        -- read
			Keyboard_avalon_ps2_slave_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Keyboard_avalon_ps2_slave_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			Keyboard_avalon_ps2_slave_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			Keyboard_avalon_ps2_slave_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			Keyboard_avalon_ps2_slave_chipselect            : out std_logic;                                        -- chipselect
			LEDs_s1_address                                 : out std_logic_vector(2 downto 0);                     -- address
			LEDs_s1_write                                   : out std_logic;                                        -- write
			LEDs_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			LEDs_s1_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			LEDs_s1_chipselect                              : out std_logic;                                        -- chipselect
			Performance_Counter_control_slave_address       : out std_logic_vector(3 downto 0);                     -- address
			Performance_Counter_control_slave_write         : out std_logic;                                        -- write
			Performance_Counter_control_slave_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Performance_Counter_control_slave_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			Performance_Counter_control_slave_begintransfer : out std_logic;                                        -- begintransfer
			PLL_pll_slave_address                           : out std_logic_vector(1 downto 0);                     -- address
			PLL_pll_slave_write                             : out std_logic;                                        -- write
			PLL_pll_slave_read                              : out std_logic;                                        -- read
			PLL_pll_slave_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			PLL_pll_slave_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			Push_Button_s1_address                          : out std_logic_vector(1 downto 0);                     -- address
			Push_Button_s1_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			RAM_s1_address                                  : out std_logic_vector(9 downto 0);                     -- address
			RAM_s1_write                                    : out std_logic;                                        -- write
			RAM_s1_readdata                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			RAM_s1_writedata                                : out std_logic_vector(31 downto 0);                    -- writedata
			RAM_s1_byteenable                               : out std_logic_vector(3 downto 0);                     -- byteenable
			RAM_s1_chipselect                               : out std_logic;                                        -- chipselect
			RAM_s1_clken                                    : out std_logic;                                        -- clken
			ROM_s1_address                                  : out std_logic_vector(11 downto 0);                    -- address
			ROM_s1_write                                    : out std_logic;                                        -- write
			ROM_s1_readdata                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ROM_s1_writedata                                : out std_logic_vector(31 downto 0);                    -- writedata
			ROM_s1_byteenable                               : out std_logic_vector(3 downto 0);                     -- byteenable
			ROM_s1_chipselect                               : out std_logic;                                        -- chipselect
			ROM_s1_clken                                    : out std_logic;                                        -- clken
			ROM_s1_debugaccess                              : out std_logic;                                        -- debugaccess
			SDRAM_s1_address                                : out std_logic_vector(23 downto 0);                    -- address
			SDRAM_s1_write                                  : out std_logic;                                        -- write
			SDRAM_s1_read                                   : out std_logic;                                        -- read
			SDRAM_s1_readdata                               : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			SDRAM_s1_writedata                              : out std_logic_vector(15 downto 0);                    -- writedata
			SDRAM_s1_byteenable                             : out std_logic_vector(1 downto 0);                     -- byteenable
			SDRAM_s1_readdatavalid                          : in  std_logic                     := 'X';             -- readdatavalid
			SDRAM_s1_waitrequest                            : in  std_logic                     := 'X';             -- waitrequest
			SDRAM_s1_chipselect                             : out std_logic;                                        -- chipselect
			Timer_s1_address                                : out std_logic_vector(2 downto 0);                     -- address
			Timer_s1_write                                  : out std_logic;                                        -- write
			Timer_s1_readdata                               : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			Timer_s1_writedata                              : out std_logic_vector(15 downto 0);                    -- writedata
			Timer_s1_chipselect                             : out std_logic;                                        -- chipselect
			VGA_char_buffer_control_slave_address           : out std_logic_vector(0 downto 0);                     -- address
			VGA_char_buffer_control_slave_write             : out std_logic;                                        -- write
			VGA_char_buffer_control_slave_read              : out std_logic;                                        -- read
			VGA_char_buffer_control_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			VGA_char_buffer_control_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			VGA_char_buffer_control_slave_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			VGA_char_buffer_control_slave_chipselect        : out std_logic;                                        -- chipselect
			VGA_char_buffersource_slave_address             : out std_logic_vector(12 downto 0);                    -- address
			VGA_char_buffersource_slave_write               : out std_logic;                                        -- write
			VGA_char_buffersource_slave_read                : out std_logic;                                        -- read
			VGA_char_buffersource_slave_readdata            : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			VGA_char_buffersource_slave_writedata           : out std_logic_vector(7 downto 0);                     -- writedata
			VGA_char_buffersource_slave_byteenable          : out std_logic_vector(0 downto 0);                     -- byteenable
			VGA_char_buffersource_slave_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			VGA_char_buffersource_slave_chipselect          : out std_logic;                                        -- chipselect
			VGA_pixel_buffer_slave_address                  : out std_logic_vector(1 downto 0);                     -- address
			VGA_pixel_buffer_slave_write                    : out std_logic;                                        -- write
			VGA_pixel_buffer_slave_read                     : out std_logic;                                        -- read
			VGA_pixel_buffer_slave_readdata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			VGA_pixel_buffer_slave_writedata                : out std_logic_vector(31 downto 0);                    -- writedata
			VGA_pixel_buffer_slave_byteenable               : out std_logic_vector(3 downto 0);                     -- byteenable
			VGA_rgb_resampler_slave_read                    : out std_logic;                                        -- read
			VGA_rgb_resampler_slave_readdata                : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component EV19_SoC_mm_interconnect_0;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal pll_c0_clk                                                        : std_logic;                     -- PLL:c0 -> [ADC:clock, Dip_Switch:clk, EV19_Core_0:clock, ID:clock, Keyboard:clk, LEDs:clk, PLL:clk, Performance_Counter:clk, Push_Button:clk, RAM:clk, ROM:clk, SDRAM:clk, Timer:clk, VGA:sys_clk_clk, mm_interconnect_0:PLL_c0_clk, rst_controller:clk]
	signal pll_c2_clk                                                        : std_logic;                     -- PLL:c2 -> VGA:vga_clk_clk
	signal ev19_core_0_data_master_readdata                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:EV19_Core_0_Data_Master_readdata -> EV19_Core_0:dataMemReadData
	signal ev19_core_0_data_master_waitrequest                               : std_logic;                     -- mm_interconnect_0:EV19_Core_0_Data_Master_waitrequest -> EV19_Core_0:dataMemWaitReq
	signal ev19_core_0_data_master_address                                   : std_logic_vector(31 downto 0); -- EV19_Core_0:dataMemAddress -> mm_interconnect_0:EV19_Core_0_Data_Master_address
	signal ev19_core_0_data_master_byteenable                                : std_logic_vector(3 downto 0);  -- EV19_Core_0:dataMemByteEnable -> mm_interconnect_0:EV19_Core_0_Data_Master_byteenable
	signal ev19_core_0_data_master_read                                      : std_logic;                     -- EV19_Core_0:dataMemReadReq -> mm_interconnect_0:EV19_Core_0_Data_Master_read
	signal ev19_core_0_data_master_writedata                                 : std_logic_vector(31 downto 0); -- EV19_Core_0:dataMemWriteData -> mm_interconnect_0:EV19_Core_0_Data_Master_writedata
	signal ev19_core_0_data_master_write                                     : std_logic;                     -- EV19_Core_0:dataMemWriteReq -> mm_interconnect_0:EV19_Core_0_Data_Master_write
	signal vga_pixel_buffer_master_waitrequest                               : std_logic;                     -- mm_interconnect_0:VGA_pixel_buffer_master_waitrequest -> VGA:pixel_buffer_master_waitrequest
	signal vga_pixel_buffer_master_readdata                                  : std_logic_vector(15 downto 0); -- mm_interconnect_0:VGA_pixel_buffer_master_readdata -> VGA:pixel_buffer_master_readdata
	signal vga_pixel_buffer_master_address                                   : std_logic_vector(31 downto 0); -- VGA:pixel_buffer_master_address -> mm_interconnect_0:VGA_pixel_buffer_master_address
	signal vga_pixel_buffer_master_read                                      : std_logic;                     -- VGA:pixel_buffer_master_read -> mm_interconnect_0:VGA_pixel_buffer_master_read
	signal vga_pixel_buffer_master_readdatavalid                             : std_logic;                     -- mm_interconnect_0:VGA_pixel_buffer_master_readdatavalid -> VGA:pixel_buffer_master_readdatavalid
	signal vga_pixel_buffer_master_lock                                      : std_logic;                     -- VGA:pixel_buffer_master_lock -> mm_interconnect_0:VGA_pixel_buffer_master_lock
	signal ev19_core_0_instruction_master_waitrequest                        : std_logic;                     -- mm_interconnect_0:EV19_Core_0_Instruction_Master_waitrequest -> EV19_Core_0:instMemWaitReq
	signal ev19_core_0_instruction_master_readdata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:EV19_Core_0_Instruction_Master_readdata -> EV19_Core_0:instMemReadData
	signal ev19_core_0_instruction_master_read                               : std_logic;                     -- EV19_Core_0:instMemReadReq -> mm_interconnect_0:EV19_Core_0_Instruction_Master_read
	signal ev19_core_0_instruction_master_byteenable                         : std_logic_vector(3 downto 0);  -- EV19_Core_0:instMemByteEnable -> mm_interconnect_0:EV19_Core_0_Instruction_Master_byteenable
	signal ev19_core_0_instruction_master_address                            : std_logic_vector(31 downto 0); -- EV19_Core_0:instMemAddress -> mm_interconnect_0:EV19_Core_0_Instruction_Master_address
	signal mm_interconnect_0_adc_adc_slave_readdata                          : std_logic_vector(31 downto 0); -- ADC:readdata -> mm_interconnect_0:ADC_adc_slave_readdata
	signal mm_interconnect_0_adc_adc_slave_waitrequest                       : std_logic;                     -- ADC:waitrequest -> mm_interconnect_0:ADC_adc_slave_waitrequest
	signal mm_interconnect_0_adc_adc_slave_address                           : std_logic_vector(2 downto 0);  -- mm_interconnect_0:ADC_adc_slave_address -> ADC:address
	signal mm_interconnect_0_adc_adc_slave_read                              : std_logic;                     -- mm_interconnect_0:ADC_adc_slave_read -> ADC:read
	signal mm_interconnect_0_adc_adc_slave_write                             : std_logic;                     -- mm_interconnect_0:ADC_adc_slave_write -> ADC:write
	signal mm_interconnect_0_adc_adc_slave_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:ADC_adc_slave_writedata -> ADC:writedata
	signal mm_interconnect_0_keyboard_avalon_ps2_slave_chipselect            : std_logic;                     -- mm_interconnect_0:Keyboard_avalon_ps2_slave_chipselect -> Keyboard:chipselect
	signal mm_interconnect_0_keyboard_avalon_ps2_slave_readdata              : std_logic_vector(31 downto 0); -- Keyboard:readdata -> mm_interconnect_0:Keyboard_avalon_ps2_slave_readdata
	signal mm_interconnect_0_keyboard_avalon_ps2_slave_waitrequest           : std_logic;                     -- Keyboard:waitrequest -> mm_interconnect_0:Keyboard_avalon_ps2_slave_waitrequest
	signal mm_interconnect_0_keyboard_avalon_ps2_slave_address               : std_logic_vector(0 downto 0);  -- mm_interconnect_0:Keyboard_avalon_ps2_slave_address -> Keyboard:address
	signal mm_interconnect_0_keyboard_avalon_ps2_slave_read                  : std_logic;                     -- mm_interconnect_0:Keyboard_avalon_ps2_slave_read -> Keyboard:read
	signal mm_interconnect_0_keyboard_avalon_ps2_slave_byteenable            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Keyboard_avalon_ps2_slave_byteenable -> Keyboard:byteenable
	signal mm_interconnect_0_keyboard_avalon_ps2_slave_write                 : std_logic;                     -- mm_interconnect_0:Keyboard_avalon_ps2_slave_write -> Keyboard:write
	signal mm_interconnect_0_keyboard_avalon_ps2_slave_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:Keyboard_avalon_ps2_slave_writedata -> Keyboard:writedata
	signal mm_interconnect_0_vga_char_buffer_control_slave_chipselect        : std_logic;                     -- mm_interconnect_0:VGA_char_buffer_control_slave_chipselect -> VGA:char_buffer_control_slave_chipselect
	signal mm_interconnect_0_vga_char_buffer_control_slave_readdata          : std_logic_vector(31 downto 0); -- VGA:char_buffer_control_slave_readdata -> mm_interconnect_0:VGA_char_buffer_control_slave_readdata
	signal mm_interconnect_0_vga_char_buffer_control_slave_address           : std_logic_vector(0 downto 0);  -- mm_interconnect_0:VGA_char_buffer_control_slave_address -> VGA:char_buffer_control_slave_address
	signal mm_interconnect_0_vga_char_buffer_control_slave_read              : std_logic;                     -- mm_interconnect_0:VGA_char_buffer_control_slave_read -> VGA:char_buffer_control_slave_read
	signal mm_interconnect_0_vga_char_buffer_control_slave_byteenable        : std_logic_vector(3 downto 0);  -- mm_interconnect_0:VGA_char_buffer_control_slave_byteenable -> VGA:char_buffer_control_slave_byteenable
	signal mm_interconnect_0_vga_char_buffer_control_slave_write             : std_logic;                     -- mm_interconnect_0:VGA_char_buffer_control_slave_write -> VGA:char_buffer_control_slave_write
	signal mm_interconnect_0_vga_char_buffer_control_slave_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:VGA_char_buffer_control_slave_writedata -> VGA:char_buffer_control_slave_writedata
	signal mm_interconnect_0_vga_char_buffersource_slave_chipselect          : std_logic;                     -- mm_interconnect_0:VGA_char_buffersource_slave_chipselect -> VGA:char_buffersource_slave_chipselect
	signal mm_interconnect_0_vga_char_buffersource_slave_readdata            : std_logic_vector(7 downto 0);  -- VGA:char_buffersource_slave_readdata -> mm_interconnect_0:VGA_char_buffersource_slave_readdata
	signal mm_interconnect_0_vga_char_buffersource_slave_waitrequest         : std_logic;                     -- VGA:char_buffersource_slave_waitrequest -> mm_interconnect_0:VGA_char_buffersource_slave_waitrequest
	signal mm_interconnect_0_vga_char_buffersource_slave_address             : std_logic_vector(12 downto 0); -- mm_interconnect_0:VGA_char_buffersource_slave_address -> VGA:char_buffersource_slave_address
	signal mm_interconnect_0_vga_char_buffersource_slave_read                : std_logic;                     -- mm_interconnect_0:VGA_char_buffersource_slave_read -> VGA:char_buffersource_slave_read
	signal mm_interconnect_0_vga_char_buffersource_slave_byteenable          : std_logic_vector(0 downto 0);  -- mm_interconnect_0:VGA_char_buffersource_slave_byteenable -> VGA:char_buffersource_slave_byteenable
	signal mm_interconnect_0_vga_char_buffersource_slave_write               : std_logic;                     -- mm_interconnect_0:VGA_char_buffersource_slave_write -> VGA:char_buffersource_slave_write
	signal mm_interconnect_0_vga_char_buffersource_slave_writedata           : std_logic_vector(7 downto 0);  -- mm_interconnect_0:VGA_char_buffersource_slave_writedata -> VGA:char_buffersource_slave_writedata
	signal mm_interconnect_0_id_control_slave_readdata                       : std_logic_vector(31 downto 0); -- ID:readdata -> mm_interconnect_0:ID_control_slave_readdata
	signal mm_interconnect_0_id_control_slave_address                        : std_logic_vector(0 downto 0);  -- mm_interconnect_0:ID_control_slave_address -> ID:address
	signal mm_interconnect_0_performance_counter_control_slave_readdata      : std_logic_vector(31 downto 0); -- Performance_Counter:readdata -> mm_interconnect_0:Performance_Counter_control_slave_readdata
	signal mm_interconnect_0_performance_counter_control_slave_address       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Performance_Counter_control_slave_address -> Performance_Counter:address
	signal mm_interconnect_0_performance_counter_control_slave_begintransfer : std_logic;                     -- mm_interconnect_0:Performance_Counter_control_slave_begintransfer -> Performance_Counter:begintransfer
	signal mm_interconnect_0_performance_counter_control_slave_write         : std_logic;                     -- mm_interconnect_0:Performance_Counter_control_slave_write -> Performance_Counter:write
	signal mm_interconnect_0_performance_counter_control_slave_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_0:Performance_Counter_control_slave_writedata -> Performance_Counter:writedata
	signal mm_interconnect_0_vga_pixel_buffer_slave_readdata                 : std_logic_vector(31 downto 0); -- VGA:pixel_buffer_slave_readdata -> mm_interconnect_0:VGA_pixel_buffer_slave_readdata
	signal mm_interconnect_0_vga_pixel_buffer_slave_address                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:VGA_pixel_buffer_slave_address -> VGA:pixel_buffer_slave_address
	signal mm_interconnect_0_vga_pixel_buffer_slave_read                     : std_logic;                     -- mm_interconnect_0:VGA_pixel_buffer_slave_read -> VGA:pixel_buffer_slave_read
	signal mm_interconnect_0_vga_pixel_buffer_slave_byteenable               : std_logic_vector(3 downto 0);  -- mm_interconnect_0:VGA_pixel_buffer_slave_byteenable -> VGA:pixel_buffer_slave_byteenable
	signal mm_interconnect_0_vga_pixel_buffer_slave_write                    : std_logic;                     -- mm_interconnect_0:VGA_pixel_buffer_slave_write -> VGA:pixel_buffer_slave_write
	signal mm_interconnect_0_vga_pixel_buffer_slave_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_0:VGA_pixel_buffer_slave_writedata -> VGA:pixel_buffer_slave_writedata
	signal mm_interconnect_0_pll_pll_slave_readdata                          : std_logic_vector(31 downto 0); -- PLL:readdata -> mm_interconnect_0:PLL_pll_slave_readdata
	signal mm_interconnect_0_pll_pll_slave_address                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:PLL_pll_slave_address -> PLL:address
	signal mm_interconnect_0_pll_pll_slave_read                              : std_logic;                     -- mm_interconnect_0:PLL_pll_slave_read -> PLL:read
	signal mm_interconnect_0_pll_pll_slave_write                             : std_logic;                     -- mm_interconnect_0:PLL_pll_slave_write -> PLL:write
	signal mm_interconnect_0_pll_pll_slave_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:PLL_pll_slave_writedata -> PLL:writedata
	signal mm_interconnect_0_vga_rgb_resampler_slave_readdata                : std_logic_vector(31 downto 0); -- VGA:rgb_resampler_slave_readdata -> mm_interconnect_0:VGA_rgb_resampler_slave_readdata
	signal mm_interconnect_0_vga_rgb_resampler_slave_read                    : std_logic;                     -- mm_interconnect_0:VGA_rgb_resampler_slave_read -> VGA:rgb_resampler_slave_read
	signal mm_interconnect_0_leds_s1_chipselect                              : std_logic;                     -- mm_interconnect_0:LEDs_s1_chipselect -> LEDs:chipselect
	signal mm_interconnect_0_leds_s1_readdata                                : std_logic_vector(31 downto 0); -- LEDs:readdata -> mm_interconnect_0:LEDs_s1_readdata
	signal mm_interconnect_0_leds_s1_address                                 : std_logic_vector(2 downto 0);  -- mm_interconnect_0:LEDs_s1_address -> LEDs:address
	signal mm_interconnect_0_leds_s1_write                                   : std_logic;                     -- mm_interconnect_0:LEDs_s1_write -> mm_interconnect_0_leds_s1_write:in
	signal mm_interconnect_0_leds_s1_writedata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:LEDs_s1_writedata -> LEDs:writedata
	signal mm_interconnect_0_dip_switch_s1_readdata                          : std_logic_vector(31 downto 0); -- Dip_Switch:readdata -> mm_interconnect_0:Dip_Switch_s1_readdata
	signal mm_interconnect_0_dip_switch_s1_address                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Dip_Switch_s1_address -> Dip_Switch:address
	signal mm_interconnect_0_push_button_s1_readdata                         : std_logic_vector(31 downto 0); -- Push_Button:readdata -> mm_interconnect_0:Push_Button_s1_readdata
	signal mm_interconnect_0_push_button_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Push_Button_s1_address -> Push_Button:address
	signal mm_interconnect_0_timer_s1_chipselect                             : std_logic;                     -- mm_interconnect_0:Timer_s1_chipselect -> Timer:chipselect
	signal mm_interconnect_0_timer_s1_readdata                               : std_logic_vector(15 downto 0); -- Timer:readdata -> mm_interconnect_0:Timer_s1_readdata
	signal mm_interconnect_0_timer_s1_address                                : std_logic_vector(2 downto 0);  -- mm_interconnect_0:Timer_s1_address -> Timer:address
	signal mm_interconnect_0_timer_s1_write                                  : std_logic;                     -- mm_interconnect_0:Timer_s1_write -> mm_interconnect_0_timer_s1_write:in
	signal mm_interconnect_0_timer_s1_writedata                              : std_logic_vector(15 downto 0); -- mm_interconnect_0:Timer_s1_writedata -> Timer:writedata
	signal mm_interconnect_0_rom_s1_chipselect                               : std_logic;                     -- mm_interconnect_0:ROM_s1_chipselect -> ROM:chipselect
	signal mm_interconnect_0_rom_s1_readdata                                 : std_logic_vector(31 downto 0); -- ROM:readdata -> mm_interconnect_0:ROM_s1_readdata
	signal mm_interconnect_0_rom_s1_debugaccess                              : std_logic;                     -- mm_interconnect_0:ROM_s1_debugaccess -> ROM:debugaccess
	signal mm_interconnect_0_rom_s1_address                                  : std_logic_vector(11 downto 0); -- mm_interconnect_0:ROM_s1_address -> ROM:address
	signal mm_interconnect_0_rom_s1_byteenable                               : std_logic_vector(3 downto 0);  -- mm_interconnect_0:ROM_s1_byteenable -> ROM:byteenable
	signal mm_interconnect_0_rom_s1_write                                    : std_logic;                     -- mm_interconnect_0:ROM_s1_write -> ROM:write
	signal mm_interconnect_0_rom_s1_writedata                                : std_logic_vector(31 downto 0); -- mm_interconnect_0:ROM_s1_writedata -> ROM:writedata
	signal mm_interconnect_0_rom_s1_clken                                    : std_logic;                     -- mm_interconnect_0:ROM_s1_clken -> ROM:clken
	signal mm_interconnect_0_ram_s1_chipselect                               : std_logic;                     -- mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	signal mm_interconnect_0_ram_s1_readdata                                 : std_logic_vector(31 downto 0); -- RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	signal mm_interconnect_0_ram_s1_address                                  : std_logic_vector(9 downto 0);  -- mm_interconnect_0:RAM_s1_address -> RAM:address
	signal mm_interconnect_0_ram_s1_byteenable                               : std_logic_vector(3 downto 0);  -- mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	signal mm_interconnect_0_ram_s1_write                                    : std_logic;                     -- mm_interconnect_0:RAM_s1_write -> RAM:write
	signal mm_interconnect_0_ram_s1_writedata                                : std_logic_vector(31 downto 0); -- mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	signal mm_interconnect_0_ram_s1_clken                                    : std_logic;                     -- mm_interconnect_0:RAM_s1_clken -> RAM:clken
	signal mm_interconnect_0_sdram_s1_chipselect                             : std_logic;                     -- mm_interconnect_0:SDRAM_s1_chipselect -> SDRAM:az_cs
	signal mm_interconnect_0_sdram_s1_readdata                               : std_logic_vector(15 downto 0); -- SDRAM:za_data -> mm_interconnect_0:SDRAM_s1_readdata
	signal mm_interconnect_0_sdram_s1_waitrequest                            : std_logic;                     -- SDRAM:za_waitrequest -> mm_interconnect_0:SDRAM_s1_waitrequest
	signal mm_interconnect_0_sdram_s1_address                                : std_logic_vector(23 downto 0); -- mm_interconnect_0:SDRAM_s1_address -> SDRAM:az_addr
	signal mm_interconnect_0_sdram_s1_read                                   : std_logic;                     -- mm_interconnect_0:SDRAM_s1_read -> mm_interconnect_0_sdram_s1_read:in
	signal mm_interconnect_0_sdram_s1_byteenable                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:SDRAM_s1_byteenable -> mm_interconnect_0_sdram_s1_byteenable:in
	signal mm_interconnect_0_sdram_s1_readdatavalid                          : std_logic;                     -- SDRAM:za_valid -> mm_interconnect_0:SDRAM_s1_readdatavalid
	signal mm_interconnect_0_sdram_s1_write                                  : std_logic;                     -- mm_interconnect_0:SDRAM_s1_write -> mm_interconnect_0_sdram_s1_write:in
	signal mm_interconnect_0_sdram_s1_writedata                              : std_logic_vector(15 downto 0); -- mm_interconnect_0:SDRAM_s1_writedata -> SDRAM:az_data
	signal rst_controller_reset_out_reset                                    : std_logic;                     -- rst_controller:reset_out -> [ADC:reset, EV19_Core_0:reset, Keyboard:reset, PLL:reset, RAM:reset, ROM:reset, mm_interconnect_0:EV19_Core_0_reset_reset_bridge_in_reset_reset, mm_interconnect_0:VGA_sys_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                : std_logic;                     -- rst_controller:reset_req -> [ROM:reset_req, rst_translator:reset_req_in]
	signal reset_reset_n_ports_inv                                           : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_leds_s1_write_ports_inv                         : std_logic;                     -- mm_interconnect_0_leds_s1_write:inv -> LEDs:write_n
	signal mm_interconnect_0_timer_s1_write_ports_inv                        : std_logic;                     -- mm_interconnect_0_timer_s1_write:inv -> Timer:write_n
	signal mm_interconnect_0_sdram_s1_read_ports_inv                         : std_logic;                     -- mm_interconnect_0_sdram_s1_read:inv -> SDRAM:az_rd_n
	signal mm_interconnect_0_sdram_s1_byteenable_ports_inv                   : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_s1_byteenable:inv -> SDRAM:az_be_n
	signal mm_interconnect_0_sdram_s1_write_ports_inv                        : std_logic;                     -- mm_interconnect_0_sdram_s1_write:inv -> SDRAM:az_wr_n
	signal rst_controller_reset_out_reset_ports_inv                          : std_logic;                     -- rst_controller_reset_out_reset:inv -> [Dip_Switch:reset_n, ID:reset_n, LEDs:reset_n, Performance_Counter:reset_n, Push_Button:reset_n, SDRAM:reset_n, Timer:reset_n]

begin

	adc : component EV19_SoC_ADC
		generic map (
			board          => "DE0-Nano",
			board_rev      => "Autodetect",
			tsclk          => 16,
			numch          => 8,
			max10pllmultby => 1,
			max10plldivby  => 1
		)
		port map (
			clock       => pll_c0_clk,                                  --                clk.clk
			reset       => rst_controller_reset_out_reset,              --              reset.reset
			write       => mm_interconnect_0_adc_adc_slave_write,       --          adc_slave.write
			readdata    => mm_interconnect_0_adc_adc_slave_readdata,    --                   .readdata
			writedata   => mm_interconnect_0_adc_adc_slave_writedata,   --                   .writedata
			address     => mm_interconnect_0_adc_adc_slave_address,     --                   .address
			waitrequest => mm_interconnect_0_adc_adc_slave_waitrequest, --                   .waitrequest
			read        => mm_interconnect_0_adc_adc_slave_read,        --                   .read
			adc_sclk    => adc_0_external_interface_sclk,               -- external_interface.export
			adc_cs_n    => adc_0_external_interface_cs_n,               --                   .export
			adc_dout    => adc_0_external_interface_dout,               --                   .export
			adc_din     => adc_0_external_interface_din                 --                   .export
		);

	dip_switch : component EV19_SoC_Dip_Switch
		port map (
			clk      => pll_c0_clk,                               --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_dip_switch_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_dip_switch_s1_readdata, --                    .readdata
			in_port  => dip_export                                -- external_connection.export
		);

	ev19_core_0 : component Core
		port map (
			reset             => rst_controller_reset_out_reset,             --              reset.reset
			dataMemAddress    => ev19_core_0_data_master_address,            --        Data_Master.address
			dataMemByteEnable => ev19_core_0_data_master_byteenable,         --                   .byteenable
			dataMemReadData   => ev19_core_0_data_master_readdata,           --                   .readdata
			dataMemReadReq    => ev19_core_0_data_master_read,               --                   .read
			dataMemWaitReq    => ev19_core_0_data_master_waitrequest,        --                   .waitrequest
			dataMemWriteData  => ev19_core_0_data_master_writedata,          --                   .writedata
			dataMemWriteReq   => ev19_core_0_data_master_write,              --                   .write
			instMemWaitReq    => ev19_core_0_instruction_master_waitrequest, -- Instruction_Master.waitrequest
			instMemReadData   => ev19_core_0_instruction_master_readdata,    --                   .readdata
			instMemReadReq    => ev19_core_0_instruction_master_read,        --                   .read
			instMemByteEnable => ev19_core_0_instruction_master_byteenable,  --                   .byteenable
			instMemAddress    => ev19_core_0_instruction_master_address,     --                   .address
			clock             => pll_c0_clk,                                 --              clock.clk
			enablePredictor   => enablepredictor_config                      --    enablePredictor.config
		);

	id : component EV19_SoC_ID
		port map (
			clock    => pll_c0_clk,                                    --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,      --         reset.reset_n
			readdata => mm_interconnect_0_id_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_id_control_slave_address(0)  --              .address
		);

	keyboard : component EV19_SoC_Keyboard
		port map (
			clk         => pll_c0_clk,                                              --                clk.clk
			reset       => rst_controller_reset_out_reset,                          --              reset.reset
			address     => mm_interconnect_0_keyboard_avalon_ps2_slave_address(0),  --   avalon_ps2_slave.address
			chipselect  => mm_interconnect_0_keyboard_avalon_ps2_slave_chipselect,  --                   .chipselect
			byteenable  => mm_interconnect_0_keyboard_avalon_ps2_slave_byteenable,  --                   .byteenable
			read        => mm_interconnect_0_keyboard_avalon_ps2_slave_read,        --                   .read
			write       => mm_interconnect_0_keyboard_avalon_ps2_slave_write,       --                   .write
			writedata   => mm_interconnect_0_keyboard_avalon_ps2_slave_writedata,   --                   .writedata
			readdata    => mm_interconnect_0_keyboard_avalon_ps2_slave_readdata,    --                   .readdata
			waitrequest => mm_interconnect_0_keyboard_avalon_ps2_slave_waitrequest, --                   .waitrequest
			irq         => open,                                                    --          interrupt.irq
			PS2_CLK     => keyboard_CLK,                                            -- external_interface.export
			PS2_DAT     => keyboard_DAT                                             --                   .export
		);

	leds : component EV19_SoC_LEDs
		port map (
			clk        => pll_c0_clk,                                --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_leds_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_leds_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_leds_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_leds_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_leds_s1_readdata,        --                    .readdata
			out_port   => led_export                                 -- external_connection.export
		);

	pll : component EV19_SoC_PLL
		port map (
			clk                => pll_c0_clk,                                --       inclk_interface.clk
			reset              => rst_controller_reset_out_reset,            -- inclk_interface_reset.reset
			read               => mm_interconnect_0_pll_pll_slave_read,      --             pll_slave.read
			write              => mm_interconnect_0_pll_pll_slave_write,     --                      .write
			address            => mm_interconnect_0_pll_pll_slave_address,   --                      .address
			readdata           => mm_interconnect_0_pll_pll_slave_readdata,  --                      .readdata
			writedata          => mm_interconnect_0_pll_pll_slave_writedata, --                      .writedata
			inclk0             => clk_clk,                                   --                inclk0.clk
			c0                 => pll_c0_clk,                                --                    c0.clk
			c1                 => sdram_clk_clk,                             --                    c1.clk
			c2                 => pll_c2_clk,                                --                    c2.clk
			scandone           => open,                                      --           (terminated)
			scandataout        => open,                                      --           (terminated)
			areset             => '0',                                       --           (terminated)
			locked             => open,                                      --           (terminated)
			phasedone          => open,                                      --           (terminated)
			phasecounterselect => "0000",                                    --           (terminated)
			phaseupdown        => '0',                                       --           (terminated)
			phasestep          => '0',                                       --           (terminated)
			scanclk            => '0',                                       --           (terminated)
			scanclkena         => '0',                                       --           (terminated)
			scandata           => '0',                                       --           (terminated)
			configupdate       => '0'                                        --           (terminated)
		);

	performance_counter : component EV19_SoC_Performance_Counter
		port map (
			clk           => pll_c0_clk,                                                        --           clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                          --         reset.reset_n
			address       => mm_interconnect_0_performance_counter_control_slave_address,       -- control_slave.address
			begintransfer => mm_interconnect_0_performance_counter_control_slave_begintransfer, --              .begintransfer
			readdata      => mm_interconnect_0_performance_counter_control_slave_readdata,      --              .readdata
			write         => mm_interconnect_0_performance_counter_control_slave_write,         --              .write
			writedata     => mm_interconnect_0_performance_counter_control_slave_writedata      --              .writedata
		);

	push_button : component EV19_SoC_Push_Button
		port map (
			clk      => pll_c0_clk,                                --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address  => mm_interconnect_0_push_button_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_push_button_s1_readdata, --                    .readdata
			in_port  => key_export                                 -- external_connection.export
		);

	ram : component EV19_SoC_RAM
		port map (
			clk        => pll_c0_clk,                          --   clk1.clk
			address    => mm_interconnect_0_ram_s1_address,    --     s1.address
			clken      => mm_interconnect_0_ram_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_ram_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_ram_s1_write,      --       .write
			readdata   => mm_interconnect_0_ram_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_ram_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_ram_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,      -- reset1.reset
			reset_req  => '0',                                 -- (terminated)
			freeze     => '0'                                  -- (terminated)
		);

	rom : component EV19_SoC_ROM
		port map (
			clk         => pll_c0_clk,                           --   clk1.clk
			address     => mm_interconnect_0_rom_s1_address,     --     s1.address
			debugaccess => mm_interconnect_0_rom_s1_debugaccess, --       .debugaccess
			clken       => mm_interconnect_0_rom_s1_clken,       --       .clken
			chipselect  => mm_interconnect_0_rom_s1_chipselect,  --       .chipselect
			write       => mm_interconnect_0_rom_s1_write,       --       .write
			readdata    => mm_interconnect_0_rom_s1_readdata,    --       .readdata
			writedata   => mm_interconnect_0_rom_s1_writedata,   --       .writedata
			byteenable  => mm_interconnect_0_rom_s1_byteenable,  --       .byteenable
			reset       => rst_controller_reset_out_reset,       -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req,   --       .reset_req
			freeze      => '0'                                   -- (terminated)
		);

	sdram : component EV19_SoC_SDRAM
		port map (
			clk            => pll_c0_clk,                                      --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,        -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_wire_addr,                                 --  wire.export
			zs_ba          => sdram_wire_ba,                                   --      .export
			zs_cas_n       => sdram_wire_cas_n,                                --      .export
			zs_cke         => sdram_wire_cke,                                  --      .export
			zs_cs_n        => sdram_wire_cs_n,                                 --      .export
			zs_dq          => sdram_wire_dq,                                   --      .export
			zs_dqm         => sdram_wire_dqm,                                  --      .export
			zs_ras_n       => sdram_wire_ras_n,                                --      .export
			zs_we_n        => sdram_wire_we_n                                  --      .export
		);

	timer : component EV19_SoC_Timer
		port map (
			clk        => pll_c0_clk,                                 --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   -- reset.reset_n
			address    => mm_interconnect_0_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_s1_write_ports_inv, --      .write_n
			irq        => open                                        --   irq.irq
		);

	vga : component EV19_SoC_VGA
		port map (
			char_buffer_control_slave_address    => mm_interconnect_0_vga_char_buffer_control_slave_address(0),  -- char_buffer_control_slave.address
			char_buffer_control_slave_byteenable => mm_interconnect_0_vga_char_buffer_control_slave_byteenable,  --                          .byteenable
			char_buffer_control_slave_chipselect => mm_interconnect_0_vga_char_buffer_control_slave_chipselect,  --                          .chipselect
			char_buffer_control_slave_read       => mm_interconnect_0_vga_char_buffer_control_slave_read,        --                          .read
			char_buffer_control_slave_write      => mm_interconnect_0_vga_char_buffer_control_slave_write,       --                          .write
			char_buffer_control_slave_writedata  => mm_interconnect_0_vga_char_buffer_control_slave_writedata,   --                          .writedata
			char_buffer_control_slave_readdata   => mm_interconnect_0_vga_char_buffer_control_slave_readdata,    --                          .readdata
			char_buffersource_slave_byteenable   => mm_interconnect_0_vga_char_buffersource_slave_byteenable(0), --   char_buffersource_slave.byteenable
			char_buffersource_slave_chipselect   => mm_interconnect_0_vga_char_buffersource_slave_chipselect,    --                          .chipselect
			char_buffersource_slave_read         => mm_interconnect_0_vga_char_buffersource_slave_read,          --                          .read
			char_buffersource_slave_write        => mm_interconnect_0_vga_char_buffersource_slave_write,         --                          .write
			char_buffersource_slave_writedata    => mm_interconnect_0_vga_char_buffersource_slave_writedata,     --                          .writedata
			char_buffersource_slave_readdata     => mm_interconnect_0_vga_char_buffersource_slave_readdata,      --                          .readdata
			char_buffersource_slave_waitrequest  => mm_interconnect_0_vga_char_buffersource_slave_waitrequest,   --                          .waitrequest
			char_buffersource_slave_address      => mm_interconnect_0_vga_char_buffersource_slave_address,       --                          .address
			pixel_buffer_master_readdatavalid    => vga_pixel_buffer_master_readdatavalid,                       --       pixel_buffer_master.readdatavalid
			pixel_buffer_master_waitrequest      => vga_pixel_buffer_master_waitrequest,                         --                          .waitrequest
			pixel_buffer_master_address          => vga_pixel_buffer_master_address,                             --                          .address
			pixel_buffer_master_lock             => vga_pixel_buffer_master_lock,                                --                          .lock
			pixel_buffer_master_read             => vga_pixel_buffer_master_read,                                --                          .read
			pixel_buffer_master_readdata         => vga_pixel_buffer_master_readdata,                            --                          .readdata
			pixel_buffer_slave_address           => mm_interconnect_0_vga_pixel_buffer_slave_address,            --        pixel_buffer_slave.address
			pixel_buffer_slave_byteenable        => mm_interconnect_0_vga_pixel_buffer_slave_byteenable,         --                          .byteenable
			pixel_buffer_slave_read              => mm_interconnect_0_vga_pixel_buffer_slave_read,               --                          .read
			pixel_buffer_slave_write             => mm_interconnect_0_vga_pixel_buffer_slave_write,              --                          .write
			pixel_buffer_slave_writedata         => mm_interconnect_0_vga_pixel_buffer_slave_writedata,          --                          .writedata
			pixel_buffer_slave_readdata          => mm_interconnect_0_vga_pixel_buffer_slave_readdata,           --                          .readdata
			rgb_resampler_slave_read             => mm_interconnect_0_vga_rgb_resampler_slave_read,              --       rgb_resampler_slave.read
			rgb_resampler_slave_readdata         => mm_interconnect_0_vga_rgb_resampler_slave_readdata,          --                          .readdata
			sys_clk_clk                          => pll_c0_clk,                                                  --                   sys_clk.clk
			sys_reset_reset_n                    => reset_reset_n,                                               --                 sys_reset.reset_n
			vga_CLK                              => vga_CLK,                                                     --                       vga.CLK
			vga_HS                               => vga_HS,                                                      --                          .HS
			vga_VS                               => vga_VS,                                                      --                          .VS
			vga_BLANK                            => vga_BLANK,                                                   --                          .BLANK
			vga_SYNC                             => vga_SYNC,                                                    --                          .SYNC
			vga_R                                => vga_R,                                                       --                          .R
			vga_G                                => vga_G,                                                       --                          .G
			vga_B                                => vga_B,                                                       --                          .B
			vga_clk_clk                          => pll_c2_clk,                                                  --                   vga_clk.clk
			vga_reset_reset_n                    => reset_reset_n                                                --                 vga_reset.reset_n
		);

	mm_interconnect_0 : component EV19_SoC_mm_interconnect_0
		port map (
			PLL_c0_clk                                      => pll_c0_clk,                                                        --                                  PLL_c0.clk
			EV19_Core_0_reset_reset_bridge_in_reset_reset   => rst_controller_reset_out_reset,                                    -- EV19_Core_0_reset_reset_bridge_in_reset.reset
			VGA_sys_reset_reset_bridge_in_reset_reset       => rst_controller_reset_out_reset,                                    --     VGA_sys_reset_reset_bridge_in_reset.reset
			EV19_Core_0_Data_Master_address                 => ev19_core_0_data_master_address,                                   --                 EV19_Core_0_Data_Master.address
			EV19_Core_0_Data_Master_waitrequest             => ev19_core_0_data_master_waitrequest,                               --                                        .waitrequest
			EV19_Core_0_Data_Master_byteenable              => ev19_core_0_data_master_byteenable,                                --                                        .byteenable
			EV19_Core_0_Data_Master_read                    => ev19_core_0_data_master_read,                                      --                                        .read
			EV19_Core_0_Data_Master_readdata                => ev19_core_0_data_master_readdata,                                  --                                        .readdata
			EV19_Core_0_Data_Master_write                   => ev19_core_0_data_master_write,                                     --                                        .write
			EV19_Core_0_Data_Master_writedata               => ev19_core_0_data_master_writedata,                                 --                                        .writedata
			EV19_Core_0_Instruction_Master_address          => ev19_core_0_instruction_master_address,                            --          EV19_Core_0_Instruction_Master.address
			EV19_Core_0_Instruction_Master_waitrequest      => ev19_core_0_instruction_master_waitrequest,                        --                                        .waitrequest
			EV19_Core_0_Instruction_Master_byteenable       => ev19_core_0_instruction_master_byteenable,                         --                                        .byteenable
			EV19_Core_0_Instruction_Master_read             => ev19_core_0_instruction_master_read,                               --                                        .read
			EV19_Core_0_Instruction_Master_readdata         => ev19_core_0_instruction_master_readdata,                           --                                        .readdata
			VGA_pixel_buffer_master_address                 => vga_pixel_buffer_master_address,                                   --                 VGA_pixel_buffer_master.address
			VGA_pixel_buffer_master_waitrequest             => vga_pixel_buffer_master_waitrequest,                               --                                        .waitrequest
			VGA_pixel_buffer_master_read                    => vga_pixel_buffer_master_read,                                      --                                        .read
			VGA_pixel_buffer_master_readdata                => vga_pixel_buffer_master_readdata,                                  --                                        .readdata
			VGA_pixel_buffer_master_readdatavalid           => vga_pixel_buffer_master_readdatavalid,                             --                                        .readdatavalid
			VGA_pixel_buffer_master_lock                    => vga_pixel_buffer_master_lock,                                      --                                        .lock
			ADC_adc_slave_address                           => mm_interconnect_0_adc_adc_slave_address,                           --                           ADC_adc_slave.address
			ADC_adc_slave_write                             => mm_interconnect_0_adc_adc_slave_write,                             --                                        .write
			ADC_adc_slave_read                              => mm_interconnect_0_adc_adc_slave_read,                              --                                        .read
			ADC_adc_slave_readdata                          => mm_interconnect_0_adc_adc_slave_readdata,                          --                                        .readdata
			ADC_adc_slave_writedata                         => mm_interconnect_0_adc_adc_slave_writedata,                         --                                        .writedata
			ADC_adc_slave_waitrequest                       => mm_interconnect_0_adc_adc_slave_waitrequest,                       --                                        .waitrequest
			Dip_Switch_s1_address                           => mm_interconnect_0_dip_switch_s1_address,                           --                           Dip_Switch_s1.address
			Dip_Switch_s1_readdata                          => mm_interconnect_0_dip_switch_s1_readdata,                          --                                        .readdata
			ID_control_slave_address                        => mm_interconnect_0_id_control_slave_address,                        --                        ID_control_slave.address
			ID_control_slave_readdata                       => mm_interconnect_0_id_control_slave_readdata,                       --                                        .readdata
			Keyboard_avalon_ps2_slave_address               => mm_interconnect_0_keyboard_avalon_ps2_slave_address,               --               Keyboard_avalon_ps2_slave.address
			Keyboard_avalon_ps2_slave_write                 => mm_interconnect_0_keyboard_avalon_ps2_slave_write,                 --                                        .write
			Keyboard_avalon_ps2_slave_read                  => mm_interconnect_0_keyboard_avalon_ps2_slave_read,                  --                                        .read
			Keyboard_avalon_ps2_slave_readdata              => mm_interconnect_0_keyboard_avalon_ps2_slave_readdata,              --                                        .readdata
			Keyboard_avalon_ps2_slave_writedata             => mm_interconnect_0_keyboard_avalon_ps2_slave_writedata,             --                                        .writedata
			Keyboard_avalon_ps2_slave_byteenable            => mm_interconnect_0_keyboard_avalon_ps2_slave_byteenable,            --                                        .byteenable
			Keyboard_avalon_ps2_slave_waitrequest           => mm_interconnect_0_keyboard_avalon_ps2_slave_waitrequest,           --                                        .waitrequest
			Keyboard_avalon_ps2_slave_chipselect            => mm_interconnect_0_keyboard_avalon_ps2_slave_chipselect,            --                                        .chipselect
			LEDs_s1_address                                 => mm_interconnect_0_leds_s1_address,                                 --                                 LEDs_s1.address
			LEDs_s1_write                                   => mm_interconnect_0_leds_s1_write,                                   --                                        .write
			LEDs_s1_readdata                                => mm_interconnect_0_leds_s1_readdata,                                --                                        .readdata
			LEDs_s1_writedata                               => mm_interconnect_0_leds_s1_writedata,                               --                                        .writedata
			LEDs_s1_chipselect                              => mm_interconnect_0_leds_s1_chipselect,                              --                                        .chipselect
			Performance_Counter_control_slave_address       => mm_interconnect_0_performance_counter_control_slave_address,       --       Performance_Counter_control_slave.address
			Performance_Counter_control_slave_write         => mm_interconnect_0_performance_counter_control_slave_write,         --                                        .write
			Performance_Counter_control_slave_readdata      => mm_interconnect_0_performance_counter_control_slave_readdata,      --                                        .readdata
			Performance_Counter_control_slave_writedata     => mm_interconnect_0_performance_counter_control_slave_writedata,     --                                        .writedata
			Performance_Counter_control_slave_begintransfer => mm_interconnect_0_performance_counter_control_slave_begintransfer, --                                        .begintransfer
			PLL_pll_slave_address                           => mm_interconnect_0_pll_pll_slave_address,                           --                           PLL_pll_slave.address
			PLL_pll_slave_write                             => mm_interconnect_0_pll_pll_slave_write,                             --                                        .write
			PLL_pll_slave_read                              => mm_interconnect_0_pll_pll_slave_read,                              --                                        .read
			PLL_pll_slave_readdata                          => mm_interconnect_0_pll_pll_slave_readdata,                          --                                        .readdata
			PLL_pll_slave_writedata                         => mm_interconnect_0_pll_pll_slave_writedata,                         --                                        .writedata
			Push_Button_s1_address                          => mm_interconnect_0_push_button_s1_address,                          --                          Push_Button_s1.address
			Push_Button_s1_readdata                         => mm_interconnect_0_push_button_s1_readdata,                         --                                        .readdata
			RAM_s1_address                                  => mm_interconnect_0_ram_s1_address,                                  --                                  RAM_s1.address
			RAM_s1_write                                    => mm_interconnect_0_ram_s1_write,                                    --                                        .write
			RAM_s1_readdata                                 => mm_interconnect_0_ram_s1_readdata,                                 --                                        .readdata
			RAM_s1_writedata                                => mm_interconnect_0_ram_s1_writedata,                                --                                        .writedata
			RAM_s1_byteenable                               => mm_interconnect_0_ram_s1_byteenable,                               --                                        .byteenable
			RAM_s1_chipselect                               => mm_interconnect_0_ram_s1_chipselect,                               --                                        .chipselect
			RAM_s1_clken                                    => mm_interconnect_0_ram_s1_clken,                                    --                                        .clken
			ROM_s1_address                                  => mm_interconnect_0_rom_s1_address,                                  --                                  ROM_s1.address
			ROM_s1_write                                    => mm_interconnect_0_rom_s1_write,                                    --                                        .write
			ROM_s1_readdata                                 => mm_interconnect_0_rom_s1_readdata,                                 --                                        .readdata
			ROM_s1_writedata                                => mm_interconnect_0_rom_s1_writedata,                                --                                        .writedata
			ROM_s1_byteenable                               => mm_interconnect_0_rom_s1_byteenable,                               --                                        .byteenable
			ROM_s1_chipselect                               => mm_interconnect_0_rom_s1_chipselect,                               --                                        .chipselect
			ROM_s1_clken                                    => mm_interconnect_0_rom_s1_clken,                                    --                                        .clken
			ROM_s1_debugaccess                              => mm_interconnect_0_rom_s1_debugaccess,                              --                                        .debugaccess
			SDRAM_s1_address                                => mm_interconnect_0_sdram_s1_address,                                --                                SDRAM_s1.address
			SDRAM_s1_write                                  => mm_interconnect_0_sdram_s1_write,                                  --                                        .write
			SDRAM_s1_read                                   => mm_interconnect_0_sdram_s1_read,                                   --                                        .read
			SDRAM_s1_readdata                               => mm_interconnect_0_sdram_s1_readdata,                               --                                        .readdata
			SDRAM_s1_writedata                              => mm_interconnect_0_sdram_s1_writedata,                              --                                        .writedata
			SDRAM_s1_byteenable                             => mm_interconnect_0_sdram_s1_byteenable,                             --                                        .byteenable
			SDRAM_s1_readdatavalid                          => mm_interconnect_0_sdram_s1_readdatavalid,                          --                                        .readdatavalid
			SDRAM_s1_waitrequest                            => mm_interconnect_0_sdram_s1_waitrequest,                            --                                        .waitrequest
			SDRAM_s1_chipselect                             => mm_interconnect_0_sdram_s1_chipselect,                             --                                        .chipselect
			Timer_s1_address                                => mm_interconnect_0_timer_s1_address,                                --                                Timer_s1.address
			Timer_s1_write                                  => mm_interconnect_0_timer_s1_write,                                  --                                        .write
			Timer_s1_readdata                               => mm_interconnect_0_timer_s1_readdata,                               --                                        .readdata
			Timer_s1_writedata                              => mm_interconnect_0_timer_s1_writedata,                              --                                        .writedata
			Timer_s1_chipselect                             => mm_interconnect_0_timer_s1_chipselect,                             --                                        .chipselect
			VGA_char_buffer_control_slave_address           => mm_interconnect_0_vga_char_buffer_control_slave_address,           --           VGA_char_buffer_control_slave.address
			VGA_char_buffer_control_slave_write             => mm_interconnect_0_vga_char_buffer_control_slave_write,             --                                        .write
			VGA_char_buffer_control_slave_read              => mm_interconnect_0_vga_char_buffer_control_slave_read,              --                                        .read
			VGA_char_buffer_control_slave_readdata          => mm_interconnect_0_vga_char_buffer_control_slave_readdata,          --                                        .readdata
			VGA_char_buffer_control_slave_writedata         => mm_interconnect_0_vga_char_buffer_control_slave_writedata,         --                                        .writedata
			VGA_char_buffer_control_slave_byteenable        => mm_interconnect_0_vga_char_buffer_control_slave_byteenable,        --                                        .byteenable
			VGA_char_buffer_control_slave_chipselect        => mm_interconnect_0_vga_char_buffer_control_slave_chipselect,        --                                        .chipselect
			VGA_char_buffersource_slave_address             => mm_interconnect_0_vga_char_buffersource_slave_address,             --             VGA_char_buffersource_slave.address
			VGA_char_buffersource_slave_write               => mm_interconnect_0_vga_char_buffersource_slave_write,               --                                        .write
			VGA_char_buffersource_slave_read                => mm_interconnect_0_vga_char_buffersource_slave_read,                --                                        .read
			VGA_char_buffersource_slave_readdata            => mm_interconnect_0_vga_char_buffersource_slave_readdata,            --                                        .readdata
			VGA_char_buffersource_slave_writedata           => mm_interconnect_0_vga_char_buffersource_slave_writedata,           --                                        .writedata
			VGA_char_buffersource_slave_byteenable          => mm_interconnect_0_vga_char_buffersource_slave_byteenable,          --                                        .byteenable
			VGA_char_buffersource_slave_waitrequest         => mm_interconnect_0_vga_char_buffersource_slave_waitrequest,         --                                        .waitrequest
			VGA_char_buffersource_slave_chipselect          => mm_interconnect_0_vga_char_buffersource_slave_chipselect,          --                                        .chipselect
			VGA_pixel_buffer_slave_address                  => mm_interconnect_0_vga_pixel_buffer_slave_address,                  --                  VGA_pixel_buffer_slave.address
			VGA_pixel_buffer_slave_write                    => mm_interconnect_0_vga_pixel_buffer_slave_write,                    --                                        .write
			VGA_pixel_buffer_slave_read                     => mm_interconnect_0_vga_pixel_buffer_slave_read,                     --                                        .read
			VGA_pixel_buffer_slave_readdata                 => mm_interconnect_0_vga_pixel_buffer_slave_readdata,                 --                                        .readdata
			VGA_pixel_buffer_slave_writedata                => mm_interconnect_0_vga_pixel_buffer_slave_writedata,                --                                        .writedata
			VGA_pixel_buffer_slave_byteenable               => mm_interconnect_0_vga_pixel_buffer_slave_byteenable,               --                                        .byteenable
			VGA_rgb_resampler_slave_read                    => mm_interconnect_0_vga_rgb_resampler_slave_read,                    --                 VGA_rgb_resampler_slave.read
			VGA_rgb_resampler_slave_readdata                => mm_interconnect_0_vga_rgb_resampler_slave_readdata                 --                                        .readdata
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => pll_c0_clk,                         --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_leds_s1_write_ports_inv <= not mm_interconnect_0_leds_s1_write;

	mm_interconnect_0_timer_s1_write_ports_inv <= not mm_interconnect_0_timer_s1_write;

	mm_interconnect_0_sdram_s1_read_ports_inv <= not mm_interconnect_0_sdram_s1_read;

	mm_interconnect_0_sdram_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_s1_byteenable;

	mm_interconnect_0_sdram_s1_write_ports_inv <= not mm_interconnect_0_sdram_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of EV19_SoC
